*DCSFQ-test

.param IB=800u
I1 0 1 pwl(0 0 5p 0 10p IB 20p IB 25p 0 45p 0 50p IB 60p IB 65p 0 85p 0 90p IB 100p IB 105p 0 125p 0 130p IB 140p IB 145p 0)
X1 1 2 DCSFQ

.subckt DCSFQ a q
.model jjmod jj(rtype=1, vg=2.8mV, cap=0.2673pF, r0=300, rn=16, icrit=0.1mA)
.param B0=1.0
.param Ic0=0.0001
.param IcRs=100u*3.50888
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LB=2p
.param LP=0.2p
.param B1=2.25
.param B2=2.25
.param B3=2.5
.param L1=1p
.param L2=3.9p
.param L3=0.6p
.param L4=1.1p
.param L5=4.5p
.param L6=2p
.param IB1=275u
.param IB2=175u
.param LB1=LB
.param LB2=LB
.param LP2=LP
.param LP3=LP
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
B1 2 3 12 jjmod area=B1
B2 5 6 13 jjmod area=B2
B3 7 8 14 jjmod area=B3
IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
LB1 3 4 LB1
LB2 7 9 LB2
L1 a 1 L1
L2 1 0 L2
L3 1 2 L3
L4 3 5 L4
L5 5 7 L5
L6 7 q L6
LP2 6 0 LP2
LP3 8 0 LP3
RB1 2 102 RB1
LRB1 102 3 LRB1
RB2 5 105 RB2
LRB2 105 6 LRB2
RB3 7 107 RB3
LRB3 107 8 LRB3
.ends DCSFQ

.tran 0.01p 160p 0 0.01p

.print DEVI I1
.print NODEV 2
.print p(B1.X1)
.print p(B2.X1)
.print p(B3.X1)